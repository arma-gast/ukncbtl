`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:49:32 03/30/2010 
// Design Name: 
// Module Name:    ppu-memctr 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ppu-memctr(
    input clk,
    input din,
    input dout,
    input sync,
    input wtbt,
    input halt,
    output rply,	 
	 inout [15:0] ad
    );


endmodule
